`include "Adder_Subtractor.v"

module Adder_Subtractor_tb;
    reg [63:0] In1,In2;
    reg Mode;
    wire [63:0] Sum;
    wire Overflow;

    Adder_Subtractor dut(.In1(In1),.In2(In2),.Mode(Mode),.Sum(Sum),.Overflow(Overflow));

    initial
    begin
        $dumpfile("Adder_Subtractor.vcd");
        $dumpvars(0, Adder_Subtractor_tb);

        $monitor("At Time = %2t:\n \tIn1 = %64b(%d),\n \tIn2 = %64b(%d),\n \tSum = %64b(%d),\n \tOverflow = %1b", $time, In1, In1, In2, In2, Sum, Sum, Overflow);

        // Addition:
        #2 In1 = 64'b1011011100000100100111101111110110010011010001100101111100010111; In2 = 64'b0101101111011101111011100001110101110000100100101010001100111110; Mode = 1'b0;
        #2 In1 = 64'b0100010001000101111100010100011110100100111111011100000011100010; In2 = 64'b1011110010100001100101100011100100111000111100101100110000000011; Mode = 1'b0;
        #2 In1 = 64'b1000110100101100011100110100110011001111010111010010010011011010; In2 = 64'b1110101110000100010000011011110100111110011011101010101010001101; Mode = 1'b0;
        #2 In1 = 64'b1010110100000000111001101011111110010010011111011101101011000101; In2 = 64'b0110101101101010000010000000100110101101101100000101001110010110; Mode = 1'b0;
        #2 In1 = 64'b0100001010101001000011010000111001101011101011010100111001111000; In2 = 64'b0001100011000011010100000111101001111110010001110001101100110011; Mode = 1'b0;
        #2 In1 = 64'b0110000100001001110100010111111011011101010101011010110010010000; In2 = 64'b0001110111000011111011001110111111001010010111010011101010001100; Mode = 1'b0;
        #2 In1 = 64'b0101010000000111110100100110000111111011101001100011110010111001; In2 = 64'b0111111111101000000100011100110110011100000111100001111011000010; Mode = 1'b0;
        #2 In1 = 64'b0000100100000101100011001001000110010011100000010000100010001001; In2 = 64'b0110000010001010001000111101101011100010011000000101100001010111; Mode = 1'b0;
        #2 In1 = 64'b0010001100100010010000111111000110111101111010001100101110111100; In2 = 64'b1000101100010010111101001001010111111110000110111110110010110100; Mode = 1'b0;
        #2 In1 = 64'b0010010001011010101011001000110111000111011010101111011001010001; In2 = 64'b0010000110001101110001110111010001110101110101001001001110010111; Mode = 1'b0;

        // Subtraction:
        #2 In1 = 64'b1011011100000100100111101111110110010011010001100101111100010111; In2 = 64'b0101101111011101111011100001110101110000100100101010001100111110; Mode = 1'b1;
        #2 In1 = 64'b0100010001000101111100010100011110100100111111011100000011100010; In2 = 64'b1011110010100001100101100011100100111000111100101100110000000011; Mode = 1'b1;
        #2 In1 = 64'b1000110100101100011100110100110011001111010111010010010011011010; In2 = 64'b1110101110000100010000011011110100111110011011101010101010001101; Mode = 1'b1;
        #2 In1 = 64'b1010110100000000111001101011111110010010011111011101101011000101; In2 = 64'b0110101101101010000010000000100110101101101100000101001110010110; Mode = 1'b1;
        #2 In1 = 64'b0100001010101001000011010000111001101011101011010100111001111000; In2 = 64'b0001100011000011010100000111101001111110010001110001101100110011; Mode = 1'b1;
        #2 In1 = 64'b0110000100001001110100010111111011011101010101011010110010010000; In2 = 64'b0001110111000011111011001110111111001010010111010011101010001100; Mode = 1'b1;
        #2 In1 = 64'b0101010000000111110100100110000111111011101001100011110010111001; In2 = 64'b0111111111101000000100011100110110011100000111100001111011000010; Mode = 1'b1;
        #2 In1 = 64'b0000100100000101100011001001000110010011100000010000100010001001; In2 = 64'b0110000010001010001000111101101011100010011000000101100001010111; Mode = 1'b1;
        #2 In1 = 64'b0010001100100010010000111111000110111101111010001100101110111100; In2 = 64'b1000101100010010111101001001010111111110000110111110110010110100; Mode = 1'b1;
        #2 In1 = 64'b0010010001011010101011001000110111000111011010101111011001010001; In2 = 64'b0010000110001101110001110111010001110101110101001001001110010111; Mode = 1'b1;

        #2 $finish;
    end
endmodule