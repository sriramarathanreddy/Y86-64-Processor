`include "Xor.v"

module Xor_tb;
    reg [63:0] In1,In2;
    wire [63:0] Out;

    Xor dut(.In1(In1), .In2(In2), .Out(Out),.Overflow(Overflow));

    initial
    begin
        $dumpfile("Xor.vcd");
        $dumpvars(0, Xor_tb);

        $monitor("At Time = %2t:\n \tIn1 = %64b (%d),\n \tIn2 = %64b (%d),\n \tOut = %64b (%d),\n \tOverflow = %b", $time, In1, In1, In2, In2, Out, Out, Overflow);
        
        #2 In1 = 64'b0011000101010110100110010000011100001110010001001011101000101011; In2 = 64'b0010100101001000010101111001100000100010110100110111100001010001;
        #2 In1 = 64'b1001101010110110000010111111100100011110100100011001000011111111; In2 = 64'b0100001100001110000011010011110111010011110110100101101001001100;
        #2 In1 = 64'b1011011111111011011000100100101111111010101101001011100001010110; In2 = 64'b0010101111111100000011011011111101001010101011111101010010110101;
        #2 In1 = 64'b0101111110010100100111010101011010001111010011101011110111000001; In2 = 64'b0001111100101110100111111011001101111100100100111111000110100101;
        #2 In1 = 64'b1011010111100010111011101100000011100010110010110011001010000001; In2 = 64'b1010010011000110100000000011110011100011011111011111010010111110;
        #2 In1 = 64'b0111001101001111110010100011100001101011111100010000011111100111; In2 = 64'b0111011110101101001111110001010110010010001010110111000110001000;
        #2 In1 = 64'b1101101100000101000000000010011101011010000011010000001101000000; In2 = 64'b1010101110001011011000011010010011011011000111101000100010011111;
        #2 In1 = 64'b1111110110001001111111001110011000000001111111000000100000101010; In2 = 64'b0000011110101011101000011111011111011101001001010011001011001000;
        #2 In1 = 64'b1001011111100101011101101101011100000100101000101001101011010101; In2 = 64'b1011001101101110001011011010000101010001101010110011011100001101;
        #2 In1 = 64'b1011001111000010101101100110110101110101100001011111000101001110; In2 = 64'b1001011111110010001010011001110100010101101100001101101011000011;
        #2 $finish;
    end
endmodule