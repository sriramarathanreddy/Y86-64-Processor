`include "And.v"

module And_tb;
    reg [63:0] In1,In2;
    wire [63:0] Out;

    And dut(.In1(In1), .In2(In2), .Out(Out), .Overflow(Overflow));

    initial
    begin
        $dumpfile("And.vcd");
        $dumpvars(0, And_tb);

        $monitor("At Time = %2t:\n \tIn1 = %64b(%d),\n \tIn2 = %64b(%d),\n \tOut = %64b(%d),\n \tOverflow = %b", $time, In1, In1, In2, In2, Out, Out, Overflow);
        
        #2 In1 = 64'b0110001111000011001001100000101110100001010111011110000100010010; In2 = 64'b0100100010001101111011011001011000101001000011001010110001101000;
        #2 In1 = 64'b1100100111010011011010000011100111101011111010000011000101101101; In2 = 64'b1001100000000100001101100100001110110111110011011110000111000101;
        #2 In1 = 64'b1110110011010011010011001001010010000010010010100100111001011010; In2 = 64'b1010010001110111000011101000001001001100000101111100111111001100;
        #2 In1 = 64'b1111100010100110110110010010111010100001001010101101001110001000; In2 = 64'b1011010000001101101011111110100000010101100010000001001110001100;
        #2 In1 = 64'b1000000011010010100001000011001100001010011111000101000111010111; In2 = 64'b0100100110010101000100111110111111010111110101101110101100001011;
        #2 In1 = 64'b0110010101000101001001001101100101100100110011111100000101100111; In2 = 64'b1001101110110010010100011000111101110010001101110111110111101110;
        #2 In1 = 64'b0010000000101010100010000011000001100011111111011110010000000101; In2 = 64'b1110011000000001010011011110011011011110011001101111010010110010;
        #2 In1 = 64'b0010101101000011001001000011100100001111010100001000000101110100; In2 = 64'b1011001111001110000101110111101010100101110000100001100111100001;
        #2 In1 = 64'b1011000111100100001100000001000100000001011111010011000100101010; In2 = 64'b0010110000101100001010111001001011101110101011101010010111100001;
        #2 In1 = 64'b0111110000010001100001100011111111011011000101000111110101011001; In2 = 64'b1001001010100000100010011110111100010001110100110000101010111101;

        #2 $finish;
    end
endmodule