module And (In1,In2,Out,Overflow);
    parameter N = 64;
    input [N-1:0] In1,In2;
    output [N-1:0]Out;
    output Overflow;
    
    genvar i;
    generate
        for (i = 0; i < N; i = i + 1)
            and x1(Out[i], In1[i], In2[i]);
    endgenerate
    assign Overflow = 1'b0;
endmodule